magic
tech sky130A
timestamp 1704960849
<< nwell >>
rect -90 -150 75 550
<< nmos >>
rect -15 -400 0 -200
<< pmos >>
rect -15 -100 0 400
<< ndiff >>
rect -70 -210 -15 -200
rect -70 -390 -60 -210
rect -30 -390 -15 -210
rect -70 -400 -15 -390
rect 0 -210 55 -200
rect 0 -390 15 -210
rect 45 -390 55 -210
rect 0 -400 55 -390
<< pdiff >>
rect -70 390 -15 400
rect -70 -90 -60 390
rect -30 -90 -15 390
rect -70 -100 -15 -90
rect 0 390 55 400
rect 0 -90 15 390
rect 45 -90 55 390
rect 0 -100 55 -90
<< ndiffc >>
rect -60 -390 -30 -210
rect 15 -390 45 -210
<< pdiffc >>
rect -60 -90 -30 390
rect 15 -90 45 390
<< psubdiff >>
rect -70 -455 55 -440
rect -70 -505 -55 -455
rect 40 -505 55 -455
rect -70 -520 55 -505
<< nsubdiff >>
rect -70 515 55 530
rect -70 465 -55 515
rect 40 465 55 515
rect -70 450 55 465
<< psubdiffcont >>
rect -55 -505 40 -455
<< nsubdiffcont >>
rect -55 465 40 515
<< poly >>
rect -15 400 0 420
rect -15 -120 0 -100
rect -55 -130 0 -120
rect -55 -170 -50 -130
rect -15 -170 0 -130
rect -55 -180 0 -170
rect -15 -200 0 -180
rect -15 -420 0 -400
<< polycont >>
rect -50 -170 -15 -130
<< locali >>
rect -70 515 55 530
rect -70 465 -55 515
rect 40 465 55 515
rect -70 450 55 465
rect -70 390 -20 450
rect -70 -90 -60 390
rect -30 -90 -20 390
rect -70 -100 -20 -90
rect 5 390 55 400
rect 5 -90 15 390
rect 45 -90 55 390
rect -90 -130 -15 -120
rect -90 -170 -85 -130
rect -90 -180 -15 -170
rect 5 -130 55 -90
rect 5 -170 15 -130
rect 45 -170 55 -130
rect -70 -210 -20 -200
rect -70 -390 -60 -210
rect -30 -390 -20 -210
rect -70 -440 -20 -390
rect 5 -210 55 -170
rect 5 -390 15 -210
rect 45 -390 55 -210
rect 5 -400 55 -390
rect -70 -455 55 -440
rect -70 -505 -55 -455
rect 40 -505 55 -455
rect -70 -520 55 -505
<< viali >>
rect -55 465 40 515
rect -85 -170 -50 -130
rect 15 -170 45 -130
rect -55 -505 40 -455
<< metal1 >>
rect -455 515 410 530
rect -455 465 -55 515
rect 40 465 410 515
rect -455 450 410 465
rect -395 -130 -35 -120
rect -395 -170 -85 -130
rect -50 -170 -35 -130
rect -395 -180 -35 -170
rect 5 -130 410 -120
rect 5 -170 15 -130
rect 45 -170 410 -130
rect 5 -180 410 -170
rect -455 -455 410 -440
rect -455 -505 -55 -455
rect 40 -505 410 -455
rect -455 -520 410 -505
<< labels >>
rlabel metal1 320 490 320 490 1 vdd
rlabel metal1 335 -480 335 -480 1 vss
rlabel metal1 375 -170 400 -130 1 out
rlabel metal1 -385 -170 -360 -130 1 in
<< end >>
